module vraylib

$if linux {
}

$if windows {
}

$if macos {
}
